/***************************************************************************************************************
***************************************************************************************************************/

interface spdif_ifc (input logic rstn);

	logic audio;

endinterface : spdif_ifc
