`ifndef AHBL_SLV_DEF__SVH
`define AHBL_SLV_DEF__SVH

`define __DBG__ __DBG_AHBL_SLV__

`define HCLK        m_cfg.vifc.hclk
`define HRESETN     m_cfg.vifc.hresetn
`define HBURST      m_cfg.vifc.hburst
`define HTRANS      m_cfg.vifc.htrans
`define HSIZE       m_cfg.vifc.hsize
`define HADDR       m_cfg.vifc.haddr
`define HPROT       m_cfg.vifc.hprot
`define HWDATA      m_cfg.vifc.hwdata
`define HRDATA      m_cfg.vifc.hrdata
`define HMSTLOCK    m_cfg.vifc.hmstlock
`define HREADY      m_cfg.vifc.hready
`define HRESP       m_cfg.vifc.hresp
`define HSEL        m_cfg.vifc.hsel
`define HWRITE      m_cfg.vifc.hwrite


`endif // AHBL_SLV_DEF__SVH
