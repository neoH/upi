`ifndef UPI_MDP_UDEF__SVH
`define UPI_MDP_UDEF__SVH

`undef __DBG__


`endif // UPI_MDP_UDEF__SVH
