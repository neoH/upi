`ifndef SPDIF_DEF__SVH
`define SPDIF_DEF__SVH

/************************************************************************************************
	A file for macro definition.
************************************************************************************************/


`define RESET    m_cfg.vifc.rstn
`define LINE     m_cfg.vifc.audio
`define __DBG__  __DBG_SPDIF_BIC__


`endif // SPDIF_DEF__SVH
