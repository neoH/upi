`ifndef UPI_ADP_PKG__SV
`define UPI_ADP_PKG__SV

package upi_adp_pkg;


endpackage : upi_adp_pkg

`endif // UPI_ADP_PKG__SV
