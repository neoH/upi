/****************************************************************************************************
****************************************************************************************************/


`ifndef UPI_ADP__SVH
`define UPI_ADP__SVH


class upi_adp extends uvm_agent;



endclass : upi_adp

`endif // UPI_ADP__SVH
