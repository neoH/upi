`ifndef UPI_MDP_DEF__SVH
`define UPI_MDP_DEF__SVH


`define __DBG__ __DBG_UPI_MDP__


`endif // UPI_MDP_DEF__SVH
