`ifndef UPI__SV
`define UPI__SV

// first include all bic packages, which to include the bic_pkg.sv
`include "bic/bic_pkg.sv"

`include "data/mdp/upi_mdp_pkg.sv"

`endif // UPI__SV
