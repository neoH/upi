`ifndef UPI_ADP_DEF__SVH
`define UPI_ADP_DEF__SVH


`define __DBG__ __DBG_UPI_ADP__


`endif // UPI_ADP_DEF__SVH
