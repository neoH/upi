`ifndef UPI_MDP_PKG__SV
`define UPI_MDP_PKG__SV


package upi_mdp_pkg;

	import uvm_pkg::*;
	import bic_pkg::*;

	`include "include/type.svh"

	`include "data/mdp/upi_mdp_def.svh"

	`include "data/mdp/upi_mdp_type.svh"
	`include "data/mdp/upi_mdp_cfg.svh"
	`include "data/mdp/upi_mdp.svh"


	`include "data/mdp/upi_mdp_udef.svh"


endpackage : upi_mdp_pkg

`endif // UPI_MDP_PKG__SV
