/*********************************************************************************************************
*********************************************************************************************************/



`ifndef SPDIF_DRV__SVH
`define SPDIF_DRV__SVH

class spdif_drv extends bic_driver;




endclass : spdif_drv

`endif // SPDIF_DRV__SVH
