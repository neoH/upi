
/*********************************************************************************************************
	File to undefine the local definition.
*********************************************************************************************************/

`undef RESET
`undef LINE
`undef __DBG__
