`ifndef UPI_ADP_TYPE__SVH
`define UPI_ADP_TYPE__SVH


// upi_adp_bic_enum
//
typedef enum
{
	SPDIF,
	TDM,
	IIS,
	PCM
} upi_adp_bic_enum;


`endif // UPI_ADP_TYPE__SVH
