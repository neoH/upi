`ifndef AHBL_SLV_UDEF__SVH
`define AHBL_SLV_UDEF__SVH

`undef __DBG__

`undef HCLK
`undef HRESETN
`undef HBURST
`undef HTRANS
`undef HSIZE
`undef HADDR
`undef HPROT
`undef HWDATA
`undef HRDATA
`undef HMSTLOCK
`undef HREADY
`undef HRESP
`undef HSEL
`undef HWRITE


`endif // AHBL_SLV_UDEF__SVH
